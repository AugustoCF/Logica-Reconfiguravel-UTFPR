DIV_CLK_inst : DIV_CLK PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
