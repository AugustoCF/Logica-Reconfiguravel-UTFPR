COMP_STATE_5_inst : COMP_STATE_5 PORT MAP (
		dataa	 => dataa_sig,
		aeb	 => aeb_sig
	);
