-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.


-- Generated by Quartus Prime Version 18.1 (Build Build 625 09/12/2018)
-- Created on Wed Feb 19 23:58:20 2025

Line_Robot Line_Robot_inst
(
	.clock(clock_sig) ,	// input  clock_sig
	.reset(reset_sig) ,	// input  reset_sig
	.SE(SE_sig) ,	// input  SE_sig
	.SD(SD_sig) ,	// input  SD_sig
	.ME2(ME2_sig) ,	// output  ME2_sig
	.ME1(ME1_sig) ,	// output  ME1_sig
	.MD2(MD2_sig) ,	// output  MD2_sig
	.MD1(MD1_sig) ,	// output  MD1_sig
	.STATE2(STATE2_sig) ,	// output  STATE2_sig
	.STATE1(STATE1_sig) 	// output  STATE1_sig
);

