DIV_CLK_inst : DIV_CLK PORT MAP (
		clock	 => clock_sig,
		cnt_en	 => cnt_en_sig,
		q	 => q_sig
	);
