COMP_10_SEC_inst : COMP_10_SEC PORT MAP (
		dataa	 => dataa_sig,
		aeb	 => aeb_sig
	);
