ROM_NUM_7SEG_inst : ROM_NUM_7SEG PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
