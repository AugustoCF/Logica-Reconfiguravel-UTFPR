// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// Created on Wed Feb 19 23:58:12 2025

// synthesis message_off 10175

`timescale 1ns/1ns

module Line_Robot (
    clock,reset,SE,SD,
    ME2,ME1,MD2,MD1,STATE2,STATE1);

    input clock;
    input reset;
    input SE;
    input SD;
    tri0 reset;
    tri0 SE;
    tri0 SD;
    output ME2;
    output ME1;
    output MD2;
    output MD1;
    output STATE2;
    output STATE1;
    reg ME2;
    reg ME1;
    reg MD2;
    reg MD1;
    reg STATE2;
    reg STATE1;
    reg [3:0] fstate;
    reg [3:0] reg_fstate;
    parameter STOP=0,MAX_SPEED=1,TURN_E=2,TURN_D=3;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or SE or SD)
    begin
        if (reset) begin
            reg_fstate <= STOP;
            ME2 <= 1'b0;
            ME1 <= 1'b0;
            MD2 <= 1'b0;
            MD1 <= 1'b0;
            STATE2 <= 1'b0;
            STATE1 <= 1'b0;
        end
        else begin
            ME2 <= 1'b0;
            ME1 <= 1'b0;
            MD2 <= 1'b0;
            MD1 <= 1'b0;
            STATE2 <= 1'b0;
            STATE1 <= 1'b0;
            case (fstate)
                STOP: begin
                    if ((~(SE) & ~(SD)))
                        reg_fstate <= STOP;
                    else if ((SE & SD))
                        reg_fstate <= MAX_SPEED;
                    else if ((SE & ~(SD)))
                        reg_fstate <= TURN_E;
                    else if ((~(SE) & SD))
                        reg_fstate <= TURN_D;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= STOP;

                    MD1 <= 1'b0;

                    MD2 <= 1'b0;

                    ME1 <= 1'b0;

                    ME2 <= 1'b0;

                    STATE1 <= 1'b0;

                    STATE2 <= 1'b0;
                end
                MAX_SPEED: begin
                    if ((SE & SD))
                        reg_fstate <= MAX_SPEED;
                    else if ((~(SE) & ~(SD)))
                        reg_fstate <= STOP;
                    else if ((SE & ~(SD)))
                        reg_fstate <= TURN_E;
                    else if ((~(SE) & SD))
                        reg_fstate <= TURN_D;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= MAX_SPEED;

                    MD1 <= 1'b1;

                    MD2 <= 1'b1;

                    ME1 <= 1'b1;

                    ME2 <= 1'b1;

                    STATE1 <= 1'b1;

                    STATE2 <= 1'b1;
                end
                TURN_E: begin
                    if ((SE & ~(SD)))
                        reg_fstate <= TURN_E;
                    else if ((~(SE) & ~(SD)))
                        reg_fstate <= STOP;
                    else if ((SE & SD))
                        reg_fstate <= MAX_SPEED;
                    else if ((~(SE) & SD))
                        reg_fstate <= TURN_D;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= TURN_E;

                    MD1 <= 1'b1;

                    MD2 <= 1'b1;

                    ME1 <= 1'b1;

                    ME2 <= 1'b0;

                    STATE1 <= 1'b0;

                    STATE2 <= 1'b1;
                end
                TURN_D: begin
                    if ((~(SE) & SD))
                        reg_fstate <= TURN_D;
                    else if ((~(SE) & ~(SD)))
                        reg_fstate <= STOP;
                    else if ((SE & SD))
                        reg_fstate <= MAX_SPEED;
                    else if ((SE & ~(SD)))
                        reg_fstate <= TURN_E;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= TURN_D;

                    MD1 <= 1'b1;

                    MD2 <= 1'b0;

                    ME1 <= 1'b1;

                    ME2 <= 1'b1;

                    STATE1 <= 1'b1;

                    STATE2 <= 1'b0;
                end
                default: begin
                    ME2 <= 1'bx;
                    ME1 <= 1'bx;
                    MD2 <= 1'bx;
                    MD1 <= 1'bx;
                    STATE2 <= 1'bx;
                    STATE1 <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // Line_Robot
