CONST_5_inst : CONST_5 PORT MAP (
		result	 => result_sig
	);
