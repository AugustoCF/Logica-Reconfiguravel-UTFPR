CONST10_inst : CONST10 PORT MAP (
		result	 => result_sig
	);
