contador_inst : contador PORT MAP (
		aclr	 => aclr_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
