CONST_4_inst : CONST_4 PORT MAP (
		result	 => result_sig
	);
