COMP_STATE_4_inst : COMP_STATE_4 PORT MAP (
		dataa	 => dataa_sig,
		aeb	 => aeb_sig
	);
