ROM_BCD_7SEG_inst : ROM_BCD_7SEG PORT MAP (
		address	 => address_sig,
		clock	 => clock_sig,
		q	 => q_sig
	);
